
// File: uart_tx.sv
//---------------------------------------------------------------------------------------
// uart transmit module  
//
//---------------------------------------------------------------------------------------

module uart_tx  
(
	clock, reset,
	ce_16, tx_data, new_tx_data, 
	ser_out, tx_busy
);
//---------------------------------------------------------------------------------------
// modules inputs and outputs 
input 			clock;			// global clock input 
input 			reset;			// global reset input 
input			ce_16;			// baud rate multiplyed by 16 - generated by baud module 
input	[7:0]	tx_data;		// data byte to transmit 
input			new_tx_data;	// asserted to indicate that there is a new data byte for transmission 
output			ser_out;		// serial data output 
output 			tx_busy;		// signs that transmitter is busy 

// internal wires 
wire ce_1;		// clock enable at bit rate 

// internal registers 
reg ser_out;
reg tx_busy;
reg [3:0]	count16;
reg [3:0]	bit_count;
reg [8:0]	data_buf;
//---------------------------------------------------------------------------------------
// module implementation 
// a counter to count 16 pulses of ce_16 to generate the ce_1 pulse 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		count16 <= 4'b0;
	else if (tx_busy & ce_16)
		count16 <= count16 + 4'b1;
	else if (~tx_busy)
		count16 <= 4'b0;
end 

// ce_1 pulse indicating output data bit should be updated 
assign ce_1 = (count16 == 4'b1111) & ce_16;

// tx_busy flag 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		tx_busy <= 1'b0;
	else if (~tx_busy & new_tx_data)
		tx_busy <= 1'b1;
	else if (tx_busy & (bit_count == 4'h9) & ce_1)
		tx_busy <= 1'b0;
end 

// output bit counter 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		bit_count <= 4'h0;
	else if (tx_busy & ce_1)
		bit_count <= bit_count + 4'h1;
	else if (~tx_busy) 
		bit_count <= 4'h0;
end 

// data shift register 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		data_buf <= 9'b0;
	else if (~tx_busy)
		data_buf <= {tx_data, 1'b0};
	else if (tx_busy & ce_1)
		data_buf <= {1'b1, data_buf[8:1]};
end 

// output data bit 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		ser_out <= 1'b1;
	else if (tx_busy)
		ser_out <= data_buf[0];
	else 
		ser_out <= 1'b1;
end 

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------

// File: uart_rx.sv
//---------------------------------------------------------------------------------------
// uart receive module  
//
//---------------------------------------------------------------------------------------

module uart_rx 
(
	clock, reset,
	ce_16, ser_in, 
	rx_data, new_rx_data 
);
//---------------------------------------------------------------------------------------
// modules inputs and outputs 
input 			clock;			// global clock input 
input 			reset;			// global reset input 
input			ce_16;			// baud rate multiplyed by 16 - generated by baud module 
input			ser_in;			// serial data input 
output	[7:0]	rx_data;		// data byte received 
output 			new_rx_data;	// signs that a new byte was received 

// internal wires 
wire ce_1;		// clock enable at bit rate 
wire ce_1_mid;	// clock enable at the middle of each bit - used to sample data 

// internal registers 
reg	[7:0] rx_data;
reg	new_rx_data;
reg [1:0] in_sync;
reg rx_busy; 
reg [3:0]	count16;
reg [3:0]	bit_count;
reg [7:0]	data_buf;
//---------------------------------------------------------------------------------------
// module implementation 
// input async input is sampled twice 
always @ (posedge clock or posedge reset)
begin 
	if (reset) 
		in_sync <= 2'b11;
	else 
		in_sync <= {in_sync[0], ser_in};
end 

// a counter to count 16 pulses of ce_16 to generate the ce_1 and ce_1_mid pulses.
// this counter is used to detect the start bit while the receiver is not receiving and 
// signs the sampling cycle during reception. 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		count16 <= 4'b0;
	else if (ce_16) 
	begin 
		if (rx_busy | (in_sync[1] == 1'b0))
			count16 <= count16 + 4'b1;
		else 
			count16 <= 4'b0;
	end 
end 

// ce_1 pulse indicating expected end of current bit 
assign ce_1 = (count16 == 4'b1111) & ce_16;
// ce_1_mid pulse indication the sampling clock cycle of the current data bit 
assign ce_1_mid = (count16 == 4'b0111) & ce_16;

// receiving busy flag 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		rx_busy <= 1'b0;
	else if (~rx_busy & ce_1_mid)
		rx_busy <= 1'b1;
	else if (rx_busy & (bit_count == 4'h8) & ce_1_mid) 
		rx_busy <= 1'b0;
end 

// bit counter 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		bit_count <= 4'h0;
	else if (~rx_busy) 
		bit_count <= 4'h0;
	else if (rx_busy & ce_1_mid)
		bit_count <= bit_count + 4'h1;
end 

// data buffer shift register 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		data_buf <= 8'h0;
	else if (rx_busy & ce_1_mid)
		data_buf <= {in_sync[1], data_buf[7:1]};
end 

// data output and flag 
always @ (posedge clock or posedge reset)
begin 
	if (reset) 
	begin 
		rx_data <= 8'h0;
		new_rx_data <= 1'b0;
	end 
	else if (rx_busy & (bit_count == 4'h8) & ce_1)
	begin 
		rx_data <= data_buf;
		new_rx_data <= 1'b1;
	end 
	else 
		new_rx_data <= 1'b0;
end 

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------

// File: uart_top.sv
//---------------------------------------------------------------------------------------
// uart top level module  
//
//---------------------------------------------------------------------------------------

module uart_top 
(
	// global signals 
	clock, reset,
	// uart serial signals 
	ser_in, ser_out,
	// transmit and receive internal interface signals 
	rx_data, new_rx_data, 
	tx_data, new_tx_data, tx_busy, 
	// baud rate configuration register - see baud_gen.v for details 
	baud_freq, baud_limit, 
	baud_clk 
);
//---------------------------------------------------------------------------------------
// modules inputs and outputs 
input 			clock;			// global clock input 
input 			reset;			// global reset input 
input			ser_in;			// serial data input 
output			ser_out;		// serial data output 
input	[7:0]	tx_data;		// data byte to transmit 
input			new_tx_data;	// asserted to indicate that there is a new data byte for transmission 
output 			tx_busy;		// signs that transmitter is busy 
output	[7:0]	rx_data;		// data byte received 
output 			new_rx_data;	// signs that a new byte was received 
input	[11:0]	baud_freq;	// baud rate setting registers - see header description 
input	[15:0]	baud_limit;
output			baud_clk;

// internal wires 
wire ce_16;		// clock enable at bit rate 

assign baud_clk = ce_16;
//---------------------------------------------------------------------------------------
// module implementation 
// baud rate generator module 
baud_gen baud_gen_1
(
	.clock(clock), .reset(reset), 
	.ce_16(ce_16), .baud_freq(baud_freq), .baud_limit(baud_limit)
);

// uart receiver 
uart_rx uart_rx_1 
(
	.clock(clock), .reset(reset), 
	.ce_16(ce_16), .ser_in(ser_in), 
	.rx_data(rx_data), .new_rx_data(new_rx_data) 
);

// uart transmitter 
uart_tx  uart_tx_1
(
	.clock(clock), .reset(reset), 
	.ce_16(ce_16), .tx_data(tx_data), .new_tx_data(new_tx_data), 
	.ser_out(ser_out), .tx_busy(tx_busy) 
);

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------

// File: uart_parser.sv
//---------------------------------------------------------------------------------------
// uart parser module  
//
//---------------------------------------------------------------------------------------

module uart_parser 
(
	// global signals 
	clock, reset,
	// transmit and receive internal interface signals from uart interface 
	rx_data, new_rx_data, 
	tx_data, new_tx_data, tx_busy, 
	// internal bus to register file 
	int_address, int_wr_data, int_write,
	int_rd_data, int_read, 
	int_req, int_gnt 
);
//---------------------------------------------------------------------------------------
// parameters 
parameter		AW = 8;			// address bus width parameter 

// modules inputs and outputs 
input 			clock;			// global clock input 
input 			reset;			// global reset input 
output	[7:0]	tx_data;		// data byte to transmit 
output			new_tx_data;	// asserted to indicate that there is a new data byte for
								// transmission 
input 			tx_busy;		// signs that transmitter is busy 
input	[7:0]	rx_data;		// data byte received 
input 			new_rx_data;	// signs that a new byte was received 
output	[AW-1:0] int_address;	// address bus to register file 
output	[7:0]	int_wr_data;	// write data to register file 
output			int_write;		// write control to register file 
output			int_read;		// read control to register file 
input	[7:0]	int_rd_data;	// data read from register file 
output			int_req;		// bus access request signal 
input			int_gnt;		// bus access grant signal 

// registered outputs
reg	[7:0] tx_data;
reg new_tx_data;
reg	[AW-1:0] int_address;
reg	[7:0] int_wr_data;
reg write_req, read_req, int_write, int_read;

// internal constants 
// define characters used by the parser 
`define CHAR_CR			8'h0d
`define CHAR_LF			8'h0a
`define CHAR_SPACE		8'h20
`define CHAR_TAB		8'h09
`define CHAR_COMMA		8'h2C
`define CHAR_R_UP		8'h52
`define CHAR_r_LO		8'h72
`define CHAR_W_UP		8'h57
`define CHAR_w_LO		8'h77
`define CHAR_0			8'h30
`define CHAR_1			8'h31
`define CHAR_2			8'h32
`define CHAR_3			8'h33
`define CHAR_4			8'h34
`define CHAR_5			8'h35
`define CHAR_6			8'h36
`define CHAR_7			8'h37
`define CHAR_8			8'h38
`define CHAR_9			8'h39
`define CHAR_A_UP		8'h41
`define CHAR_B_UP		8'h42
`define CHAR_C_UP		8'h43
`define CHAR_D_UP		8'h44
`define CHAR_E_UP		8'h45
`define CHAR_F_UP		8'h46
`define CHAR_a_LO		8'h61
`define CHAR_b_LO		8'h62
`define CHAR_c_LO		8'h63
`define CHAR_d_LO		8'h64
`define CHAR_e_LO		8'h65
`define CHAR_f_LO		8'h66

// main (receive) state machine states 
`define MAIN_IDLE		4'b0000
`define MAIN_WHITE1		4'b0001
`define MAIN_DATA		4'b0010
`define MAIN_WHITE2		4'b0011
`define MAIN_ADDR		4'b0100
`define MAIN_EOL		4'b0101
// binary mode extension states 
`define MAIN_BIN_CMD	4'b1000
`define MAIN_BIN_ADRH	4'b1001
`define MAIN_BIN_ADRL	4'b1010
`define MAIN_BIN_LEN    4'b1011
`define MAIN_BIN_DATA   4'b1100 

// transmit state machine 
`define TX_IDLE			3'b000
`define TX_HI_NIB		3'b001
`define TX_LO_NIB		3'b100
`define TX_CHAR_CR		3'b101
`define TX_CHAR_LF		3'b110

// binary extension mode commands - the command is indicated by bits 5:4 of the command byte 
`define BIN_CMD_NOP		2'b00
`define BIN_CMD_READ	2'b01
`define BIN_CMD_WRITE	2'b10

// internal wires and registers 
reg [3:0] main_sm;			// main state machine 
reg read_op;				// read operation flag 
reg write_op;				// write operation flag 
reg data_in_hex_range;		// indicates that the received data is in the range of hex number 
reg [7:0] data_param;		// operation data parameter 
reg [15:0] addr_param;		// operation address parameter 
reg [3:0] data_nibble;		// data nibble from received character 
reg read_done;				// internally generated read done flag 
reg read_done_s;			// sampled read done 
reg [7:0] read_data_s;		// sampled read data 
reg [3:0] tx_nibble;		// nibble value for transmission 
reg [7:0] tx_char;			// transmit byte from nibble to character conversion 
reg [2:0] tx_sm;			// transmit state machine 
reg s_tx_busy;				// sampled tx_busy for falling edge detection 
reg bin_read_op;			// binary mode read operation flag 
reg bin_write_op;			// binary mode write operation flag 
reg addr_auto_inc;			// address auto increment mode 
reg send_stat_flag;			// send status flag 
reg [7:0] bin_byte_count;	// binary mode byte counter 
wire bin_last_byte;			// last byte flag indicates that the current byte in the command is the last 
wire tx_end_p;				// transmission end pulse 

//---------------------------------------------------------------------------------------
// module implementation 
// main state machine 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		main_sm <= `MAIN_IDLE;
	else if (new_rx_data) 
	begin 
		case (main_sm)
			// wait for a read ('r') or write ('w') command 
			// binary extension - an all zeros byte enabled binary commands 
			`MAIN_IDLE:
				// check received character 
				if (rx_data == 8'h0)
					// an all zeros received byte enters binary mode 
					main_sm <= `MAIN_BIN_CMD;
				else if ((rx_data == `CHAR_r_LO) | (rx_data == `CHAR_R_UP))
					// on read wait to receive only address field 
					main_sm <= `MAIN_WHITE2;
				else if ((rx_data == `CHAR_w_LO) | (rx_data == `CHAR_W_UP))
					// on write wait to receive data and address 
					main_sm <= `MAIN_WHITE1;
				else if ((rx_data == `CHAR_CR) | (rx_data == `CHAR_LF))
					// on new line sta in idle 
					main_sm <= `MAIN_IDLE;
				else 
					// any other character wait to end of line (EOL)
					main_sm <= `MAIN_EOL;
				
			// wait for white spaces till first data nibble 
			`MAIN_WHITE1:
				// wait in this case until any white space character is received. in any 
				// valid character for data value switch to data state. a new line or carriage 
				// return should reset the state machine to idle.
				// any other character transitions the state machine to wait for EOL.
				if ((rx_data == `CHAR_SPACE) | (rx_data == `CHAR_TAB))
					main_sm <= `MAIN_WHITE1;
				else if (data_in_hex_range)
					main_sm <= `MAIN_DATA;
				else if ((rx_data == `CHAR_CR) | (rx_data == `CHAR_LF))
					main_sm <= `MAIN_IDLE;
				else 
					main_sm <= `MAIN_EOL;
					
			// receive data field 
			`MAIN_DATA:
				// wait while data in hex range. white space transition to wait white 2 state.
				// CR and LF resets the state machine. any other value cause state machine to 
				// wait til end of line.
				if (data_in_hex_range)
					main_sm <= `MAIN_DATA;
				else if ((rx_data == `CHAR_SPACE) | (rx_data == `CHAR_TAB))
					main_sm <= `MAIN_WHITE2;
				else if ((rx_data == `CHAR_CR) | (rx_data == `CHAR_LF))
					main_sm <= `MAIN_IDLE;
				else 
					main_sm <= `MAIN_EOL;
				
			// wait for white spaces till first address nibble 
			`MAIN_WHITE2:
				// similar to MAIN_WHITE1 
				if ((rx_data == `CHAR_SPACE) | (rx_data == `CHAR_TAB))
					main_sm <= `MAIN_WHITE2;
				else if (data_in_hex_range)
					main_sm <= `MAIN_ADDR;
				else if ((rx_data == `CHAR_CR) | (rx_data == `CHAR_LF))
					main_sm <= `MAIN_IDLE;
				else 
					main_sm <= `MAIN_EOL;

			// receive address field 
			`MAIN_ADDR:
				// similar to MAIN_DATA 
				if (data_in_hex_range)
					main_sm <= `MAIN_ADDR;
				else if ((rx_data == `CHAR_CR) | (rx_data == `CHAR_LF))
					main_sm <= `MAIN_IDLE;
				else 
					main_sm <= `MAIN_EOL;

			// wait to EOL 				
			`MAIN_EOL:
				// wait for CR or LF to move back to idle 
				if ((rx_data == `CHAR_CR) | (rx_data == `CHAR_LF))
					main_sm <= `MAIN_IDLE;
					
			// binary extension 
			// wait for command - one byte 
			`MAIN_BIN_CMD:
				// check if command is a NOP command 
				if (rx_data[5:4] == `BIN_CMD_NOP)
					// if NOP command then switch back to idle state 
					main_sm <= `MAIN_IDLE;
				else 
					// not a NOP command, continue receiving parameters 
					main_sm <= `MAIN_BIN_ADRH;
							
			// wait for address parameter - two bytes 
			// high address byte 
			`MAIN_BIN_ADRH:
				// switch to next state 
				main_sm <= `MAIN_BIN_ADRL;
			
			// low address byte 
			`MAIN_BIN_ADRL:
				// switch to next state 
				main_sm <= `MAIN_BIN_LEN;
			
			// wait for length parameter - one byte 
			`MAIN_BIN_LEN:
				// check if write command else command reception ended 
				if (bin_write_op)
					// wait for write data 
					main_sm <= `MAIN_BIN_DATA;
				else 
					// command reception has ended 
					main_sm <= `MAIN_IDLE;
			
			// on write commands wait for data till end of buffer as specified by length parameter 
			`MAIN_BIN_DATA:
				// if this is the last data byte then return to idle 
				if (bin_last_byte)
					main_sm <= `MAIN_IDLE;
				
			// go to idle 
			default:
				main_sm <= `MAIN_IDLE;
		endcase 
	end 
end 

// indicates that the received data is in the range of hex number 
always @ (rx_data)
begin 
	if (((rx_data >= `CHAR_0   ) && (rx_data <= `CHAR_9   )) || 
	    ((rx_data >= `CHAR_A_UP) && (rx_data <= `CHAR_F_UP)) || 
	    ((rx_data >= `CHAR_a_LO) && (rx_data <= `CHAR_f_LO)))
		data_in_hex_range <= 1'b1;
	else 
		data_in_hex_range <= 1'b0;
end 

// read operation flag 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		read_op <= 1'b0;
	else if ((main_sm == `MAIN_IDLE) && new_rx_data) 
	begin 
		// the read operation flag is set when a read command is received in idle state and cleared 
		// if any other character is received during that state.
		if ((rx_data == `CHAR_r_LO) | (rx_data == `CHAR_R_UP))
			read_op <= 1'b1;
		else 
			read_op <= 1'b0;
	end 
end 

// write operation flag 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		write_op <= 1'b0;
	else if ((main_sm == `MAIN_IDLE) & new_rx_data) 
	begin 
		// the write operation flag is set when a write command is received in idle state and cleared 
		// if any other character is received during that state.
		if ((rx_data == `CHAR_w_LO) | (rx_data == `CHAR_W_UP))
			write_op <= 1'b1;
		else 
			write_op <= 1'b0;
	end 
end 

// binary mode read operation flag 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		bin_read_op <= 1'b0;
	else if ((main_sm == `MAIN_BIN_CMD) && new_rx_data && (rx_data[5:4] == `BIN_CMD_READ))
		// read command is started on reception of a read command 
		bin_read_op <= 1'b1;
	else if (bin_read_op && tx_end_p && bin_last_byte)
		// read command ends on transmission of the last byte read 
		bin_read_op <= 1'b0;
end 

// binary mode write operation flag 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		bin_write_op <= 1'b0;
	else if ((main_sm == `MAIN_BIN_CMD) && new_rx_data && (rx_data[5:4] == `BIN_CMD_WRITE))
		// write command is started on reception of a write command 
		bin_write_op <= 1'b1;
	else if ((main_sm == `MAIN_BIN_DATA) && new_rx_data && bin_last_byte)
		bin_write_op <= 1'b0;
end 

// send status flag - used only in binary extension mode 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		send_stat_flag <= 1'b0;
	else if ((main_sm == `MAIN_BIN_CMD) && new_rx_data)
	begin 
		// check if a status byte should be sent at the end of the command 
		if (rx_data[0] == 1'b1)
			send_stat_flag <= 1'b1;
		else 
			send_stat_flag <= 1'b0;
	end 
end 

// address auto increment - used only in binary extension mode 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		addr_auto_inc <= 1'b0;
	else if ((main_sm == `MAIN_BIN_CMD) && new_rx_data)
	begin 
		// check if address should be automatically incremented or not. 
		// Note that when rx_data[1] is set, address auto increment is disabled. 
		if (rx_data[1] == 1'b0)
			addr_auto_inc <= 1'b1;
		else 
			addr_auto_inc <= 1'b0;
	end 
end 

// operation data parameter 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		data_param <= 8'h0;
	else if ((main_sm == `MAIN_WHITE1) & new_rx_data & data_in_hex_range) 
		data_param <= {4'h0, data_nibble};
	else if ((main_sm == `MAIN_DATA) & new_rx_data & data_in_hex_range) 
		data_param <= {data_param[3:0], data_nibble};
end 

// operation address parameter 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		addr_param <= 0;
	else if ((main_sm == `MAIN_WHITE2) & new_rx_data & data_in_hex_range) 
		addr_param <= {12'b0, data_nibble};
	else if ((main_sm == `MAIN_ADDR) & new_rx_data & data_in_hex_range) 
		addr_param <= {addr_param[11:0], data_nibble};
	// binary extension 
	else if (main_sm == `MAIN_BIN_ADRH)
		addr_param[15:8] <= rx_data;
	else if (main_sm == `MAIN_BIN_ADRL)
		addr_param[7:0] <= rx_data;
end 

// binary mode command byte counter is loaded with the length parameter and counts down to zero.
// NOTE: a value of zero for the length parameter indicates a command of 256 bytes.
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		bin_byte_count <= 8'b0;
	else if ((main_sm == `MAIN_BIN_LEN) && new_rx_data)
		bin_byte_count <= rx_data;
	else if ((bin_write_op && (main_sm == `MAIN_BIN_DATA) && new_rx_data) || 
			 (bin_read_op && tx_end_p))
		// byte counter is updated on every new data received in write operations and for every 
		// byte transmitted for read operations.
		bin_byte_count <= bin_byte_count - 1;
end 
// last byte in command flag 
assign bin_last_byte = (bin_byte_count == 8'h01) ? 1'b1 : 1'b0;

// internal write control and data 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
	begin 
		write_req <= 1'b0;
		int_write <= 1'b0;
		int_wr_data <= 0;
	end 
	else if (write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range)
	begin 
		write_req <= 1'b1;
		int_wr_data <= data_param;
	end 
	// binary extension mode 
	else if (bin_write_op && (main_sm == `MAIN_BIN_DATA) && new_rx_data) 
	begin 
		write_req <= 1'b1;
		int_wr_data <= rx_data;
	end 
	else if (int_gnt && write_req) 
	begin 
		// set internal bus write and clear the write request flag 
		int_write <= 1'b1;
		write_req <= 1'b0;
	end 
	else 
		int_write <= 1'b0;
end 

// internal read control 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
	begin 
		int_read <= 1'b0;
		read_req <= 1'b0;
	end 
	else if (read_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range)
		read_req <= 1'b1;
	// binary extension 
	else if (bin_read_op && (main_sm == `MAIN_BIN_LEN) && new_rx_data)
		// the first read request is issued on reception of the length byte 
		read_req <= 1'b1;
	else if (bin_read_op && tx_end_p && !bin_last_byte)
		// the next read requests are issued after the previous read value was transmitted and 
		// this is not the last byte to be read.
		read_req <= 1'b1;
	else if (int_gnt && read_req) 
	begin 
		// set internal bus read and clear the read request flag 
		int_read <= 1'b1;
		read_req <= 1'b0;
	end 
	else 
		int_read <= 1'b0;
end 

// external request signal is active on read or write request 
assign int_req = write_req | read_req;

// internal address 
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		int_address <= 0;
	else if ((main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range)
		int_address <= addr_param[AW-1:0];
	// binary extension 
	else if ((main_sm == `MAIN_BIN_LEN) && new_rx_data)
		// sample address parameter on reception of length byte 
		int_address <= addr_param[AW-1:0];
	else if (addr_auto_inc && 
			 ((bin_read_op && tx_end_p && !bin_last_byte) || 
			  (bin_write_op && int_write)))
		// address is incremented on every read or write if enabled 
		int_address <= int_address + 1;
end 

// read done flag and sampled data read 
always @ (posedge clock or posedge reset)
begin
	if (reset) begin 
		read_done <= 1'b0;
		read_done_s <= 1'b0;
		read_data_s <= 8'h0;
	end 
	else 
	begin 
		// read done flag 
		if (int_read) 
			read_done <= 1'b1;
		else 
			read_done <= 1'b0;
			
		// sampled read done 
		read_done_s <= read_done;
		
		// sampled data read 
		if (read_done)
			read_data_s <= int_rd_data;
	end 
end 

// transmit state machine and control 
always @ (posedge clock or posedge reset)
begin 
	if (reset) begin 
		tx_sm <= `TX_IDLE;
		tx_data <= 8'h0;
		new_tx_data <= 1'b0;
	end 
	else 
		case (tx_sm)
			// wait for read done indication 
			`TX_IDLE: 
				// on end of every read operation check how the data read should be transmitted 
				// according to read type: ascii or binary.
				if (read_done_s) 
					// on binary mode read transmit byte value 
					if (bin_read_op)
					begin 
						// note that there is no need to change state 
						tx_data <= read_data_s;
						new_tx_data <= 1'b1;
					end 
					else 
					begin 
						tx_sm <= `TX_HI_NIB;
						tx_data <= tx_char;
						new_tx_data <= 1'b1;
					end 
				// check if status byte should be transmitted 
				else if ((send_stat_flag && bin_read_op && tx_end_p && bin_last_byte) ||	// end of read command 
					(send_stat_flag && bin_write_op && new_rx_data && bin_last_byte) ||	// end of write command 
					((main_sm == `MAIN_BIN_CMD) && new_rx_data && (rx_data[5:4] == `BIN_CMD_NOP)))	// NOP 
				begin 
					// send status byte - currently a constant 
					tx_data <= 8'h5a;
					new_tx_data <= 1'b1;
				end 
				else 
					new_tx_data <= 1'b0;

			// wait for transmit to end 
			`TX_HI_NIB:	
				if (tx_end_p) 
				begin 
					tx_sm <= `TX_LO_NIB;
					tx_data <= tx_char;
					new_tx_data <= 1'b1;
				end 
				else 
					new_tx_data <= 1'b0;
					
			// wait for transmit to end 
			`TX_LO_NIB:	
				if (tx_end_p) 
				begin 
					tx_sm <= `TX_CHAR_CR;
					tx_data <= `CHAR_CR;
					new_tx_data <= 1'b1;
				end 
				else 
					new_tx_data <= 1'b0;
					
			// wait for transmit to end 
			`TX_CHAR_CR:	
				if (tx_end_p) 
				begin 
					tx_sm <= `TX_CHAR_LF;
					tx_data <= `CHAR_LF;
					new_tx_data <= 1'b1;
				end 
				else 
					new_tx_data <= 1'b0;
					
			// wait for transmit to end 
			`TX_CHAR_LF:	
				begin 
					if (tx_end_p) 
						tx_sm <= `TX_IDLE;
					// clear tx new data flag 
					new_tx_data <= 1'b0;
				end 
					
			// return to idle 
			default:
				tx_sm <= `TX_IDLE;
		endcase 
end 

// select the nibble to the nibble to character conversion 
always @ (tx_sm or read_data_s)
begin 
	case (tx_sm)
		`TX_IDLE:		tx_nibble = read_data_s[7:4];
		`TX_HI_NIB:		tx_nibble = read_data_s[3:0];
		default:		tx_nibble = read_data_s[7:4];
	endcase
end 

// sampled tx_busy 
always @ (posedge clock or posedge reset)
begin 
	if (reset)
		s_tx_busy <= 1'b0;
	else 
		s_tx_busy <= tx_busy;
end 
// tx end pulse 
assign tx_end_p = ~tx_busy & s_tx_busy;

// character to nibble conversion 
always @ (rx_data)
begin 
	case (rx_data) 
		`CHAR_0:				data_nibble = 4'h0;
		`CHAR_1:				data_nibble = 4'h1;
		`CHAR_2:				data_nibble = 4'h2;
		`CHAR_3:				data_nibble = 4'h3;
		`CHAR_4:				data_nibble = 4'h4;
		`CHAR_5:				data_nibble = 4'h5;
		`CHAR_6:				data_nibble = 4'h6;
		`CHAR_7:				data_nibble = 4'h7;
		`CHAR_8:				data_nibble = 4'h8;
		`CHAR_9:				data_nibble = 4'h9;
		`CHAR_A_UP, `CHAR_a_LO:	data_nibble = 4'ha;
		`CHAR_B_UP, `CHAR_b_LO:	data_nibble = 4'hb;
		`CHAR_C_UP, `CHAR_c_LO:	data_nibble = 4'hc;
		`CHAR_D_UP, `CHAR_d_LO:	data_nibble = 4'hd;
		`CHAR_E_UP, `CHAR_e_LO:	data_nibble = 4'he;
		`CHAR_F_UP, `CHAR_f_LO:	data_nibble = 4'hf;
		default:				data_nibble = 4'hf;
	endcase 
end 

// nibble to character conversion 
always @ (tx_nibble)
begin 
	case (tx_nibble)
		4'h0:	tx_char = `CHAR_0;
		4'h1:	tx_char = `CHAR_1;
		4'h2:	tx_char = `CHAR_2;
		4'h3:	tx_char = `CHAR_3;
		4'h4:	tx_char = `CHAR_4;
		4'h5:	tx_char = `CHAR_5;
		4'h6:	tx_char = `CHAR_6;
		4'h7:	tx_char = `CHAR_7;
		4'h8:	tx_char = `CHAR_8;
		4'h9:	tx_char = `CHAR_9;
		4'ha:	tx_char = `CHAR_A_UP;
		4'hb:	tx_char = `CHAR_B_UP;
		4'hc:	tx_char = `CHAR_C_UP;
		4'hd:	tx_char = `CHAR_D_UP;
		4'he:	tx_char = `CHAR_E_UP;
		default: tx_char = `CHAR_F_UP;
	endcase 
end 

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------

// File: uart2bus_top.sv
//---------------------------------------------------------------------------------------
// uart to internal bus top module 
//
//---------------------------------------------------------------------------------------

module uart2bus_top (
	// global signals 
	clock, reset,
	// uart serial signals 
	ser_in, ser_out,
	// internal bus to register file 
	int_address, int_wr_data, int_write,
	int_rd_data, int_read, 
	int_req, int_gnt 
);
//---------------------------------------------------------------------------------------
// modules inputs and outputs 
input 			clock;			// global clock input 
input 			reset;			// global reset input 
input			ser_in;			// serial data input 
output			ser_out;		// serial data output 
output	[15:0]	int_address;	// address bus to register file 
output	[7:0]	int_wr_data;	// write data to register file 
output			int_write;		// write control to register file 
output			int_read;		// read control to register file 
input	[7:0]	int_rd_data;	// data read from register file 
output			int_req;		// bus access request signal 
input			int_gnt;		// bus access grant signal 

// baud rate configuration, see baud_gen.v for more details.
// baud rate generator parameters for 115200 baud on 40MHz clock 
`define D_BAUD_FREQ			12'h90
`define D_BAUD_LIMIT		16'h0ba5
// baud rate generator parameters for 115200 baud on 44MHz clock 
// `define D_BAUD_FREQ			12'd23
// `define D_BAUD_LIMIT		16'd527
// baud rate generator parameters for 9600 baud on 66MHz clock 
//`define D_BAUD_FREQ		12'h10
//`define D_BAUD_LIMIT		16'h1ACB

// internal wires 
wire	[7:0]	tx_data;		// data byte to transmit 
wire			new_tx_data;	// asserted to indicate that there is a new data byte for transmission 
wire 			tx_busy;		// signs that transmitter is busy 
wire	[7:0]	rx_data;		// data byte received 
wire 			new_rx_data;	// signs that a new byte was received 
wire	[11:0]	baud_freq;
wire	[15:0]	baud_limit;
wire			baud_clk;

//---------------------------------------------------------------------------------------
// module implementation 
// uart top module instance 
uart_top uart1
(
	.clock(clock), .reset(reset),
	.ser_in(ser_in), .ser_out(ser_out),
	.rx_data(rx_data), .new_rx_data(new_rx_data), 
	.tx_data(tx_data), .new_tx_data(new_tx_data), .tx_busy(tx_busy), 
	.baud_freq(baud_freq), .baud_limit(baud_limit),
	.baud_clk(baud_clk) 
);

// assign baud rate default values 
assign baud_freq = `D_BAUD_FREQ;
assign baud_limit = `D_BAUD_LIMIT;

// uart parser instance 
uart_parser #(16) uart_parser1
(
	.clock(clock), .reset(reset),
	.rx_data(rx_data), .new_rx_data(new_rx_data), 
	.tx_data(tx_data), .new_tx_data(new_tx_data), .tx_busy(tx_busy), 
	.int_address(int_address), .int_wr_data(int_wr_data), .int_write(int_write),
	.int_rd_data(int_rd_data), .int_read(int_read), 
	.int_req(int_req), .int_gnt(int_gnt) 
);

assert_a0: assert property(@(posedge clock) int_write |-> $stable(int_wr_data));
assert_a1: assert property(@(posedge clock) $rose(int_write) |=> $stable(int_address)[*2]);
assert_a2: assert property(@(posedge clock) $rose(int_gnt) |-> ##[1:5] $fell(int_req));
assert_a3: assert property(@(posedge clock) tx_busy |-> $changed(ser_out) throughout (1'b1)[*1]);
assert_a4: assert property(@(posedge clock) $rose(int_req) |-> ##[1:2] $rose(int_gnt));
assert_a5: assert property(@(posedge clock) $rose(int_write) |=> $fell(int_write));
assert_a6: assert property(@(posedge clock) $fell(reset) |-> ##[1:5] $stable(ser_out));
assert_a7: assert property(@(posedge clock) $rose(int_read) |=> !$isunknown(int_rd_data));
assert_a8: assert property(@(posedge clock) reset |=> (ser_out == 0 && int_address == 0 && int_wr_data == 0 && int_write == 0 && int_read == 0));
assert_a9: assert property(@(posedge clock) disable iff (reset) $changed(ser_in) |-> ser_in == $past(ser_in));
assert_a10: assert property(@(posedge clock) int_write |-> ##1 !int_write);
assert_a11: assert property(@(posedge clock) int_read |-> ##1 !int_read);
assert_a12: assert property(@(posedge clock) $rose(int_read) |-> ##[1:3] $stable(int_rd_data));
assert_a13: assert property(@(posedge clock) reset |-> ser_out == 0 [*2] ##1 ser_out == 0);
assert_a14: assert property(@(posedge clock) $rose(ser_in) |-> ##[1:3] $stable(int_rd_data));
assert_a15: assert property(@(posedge clock) $fell(tx_busy) |-> ser_out ##1 ser_out ##1 ser_out);
assert_a16: assert property(@(posedge clock) $rose(int_write) |-> $past(int_wr_data, 1) == int_wr_data ##1 $future(int_wr_data, 1) == int_wr_data);
assert_a17: assert property(@(posedge clock) $changed(int_req) |-> $past(int_req) == int_req);
assert_a18: assert property(@(posedge clock) $rose(int_req) |-> $stable(int_address)[*2]);
assert_a19: assert property(@(posedge clock) $rose(int_read) |=> $fell(int_read));
assert_a20: assert property(@(posedge clock) $rose(int_req) |-> ##[1:4] $rose(int_gnt));
assert_a21: assert property(@(posedge clock) ($rose(int_write) || $rose(int_read)) |=> $stable(int_address));
assert_a22: assert property(@(posedge clock) tx_busy |-> $stable(ser_out) or $rose(ser_out) or $fell(ser_out));
assert_a23: assert property(@(posedge clock) $rose(int_write) |=> $stable(int_wr_data));
assert_a24: assert property(@(posedge clock) disable iff (reset) (uart_parser.main_sm == `MAIN_ADDR && !new_rx_data) |=> $stable(int_address));
assert_a25: assert property(@(posedge clock) $rose(!reset) |=> $stable(int_address) until_with ((uart_parser.main_sm == `MAIN_ADDR && new_rx_data && !data_in_hex_range) || (uart_parser.main_sm == `MAIN_BIN_LEN && new_rx_data) || (addr_auto_inc && ((bin_read_op && tx_end_p && !bin_last_byte) || (bin_write_op && int_write)))));
assert_a26: assert property(@(posedge clock) disable iff (reset) !( (uart_parser.main_sm == `MAIN_ADDR && new_rx_data && !data_in_hex_range) || (main_sm == `MAIN_BIN_LEN && new_rx_data) || (addr_auto_inc && ((bin_read_op && tx_end_p && !bin_last_byte) || (bin_write_op && int_write))) ) |=> $stable(int_address));
assert_a27: assert property(@(posedge clock) disable iff (reset) (addr_auto_inc && bin_read_op && tx_end_p && !bin_last_byte) |=> (int_address == $past(int_address) + 1));
assert_a28: assert property(@(posedge clock) reset |=> (int_address == 0));
assert_a29: assert property(@(posedge clock) disable iff (reset) (main_sm == `MAIN_ADDR && new_rx_data && !data_in_hex_range) |=> (int_address == $past(addr_param[AW-1:0])));
assert_a30: assert property(@(posedge clock) disable iff (reset) (main_sm == `MAIN_BIN_LEN && new_rx_data) |=> (int_address == $past(addr_param[AW-1:0])));
assert_a31: assert property(@(posedge clock) disable iff (reset) (main_sm == `MAIN_ADDR && new_rx_data && data_in_hex_range) |=> (int_address == $past(int_address)));
assert_a32: assert property(@(posedge clock) disable iff (reset) !new_rx_data |=> (int_address == $past(int_address)));
assert_a33: assert property(@(posedge clock) disable iff (reset) (bin_read_op && !addr_auto_inc && tx_end_p) |=> (int_address == $past(int_address)));
assert_a34: assert property(@(posedge clock) disable iff (reset) (addr_auto_inc && bin_write_op && int_write) |=> (int_address == $past(int_address) + 1));
assert_a35: assert property(@(posedge clock) disable iff (reset) (main_sm != `MAIN_ADDR && main_sm != `MAIN_BIN_LEN && new_rx_data) |=> (int_address == $past(int_address)));
assert_a36: assert property(@(posedge clock) disable iff (reset) ((main_sm == `MAIN_BIN_LEN) && new_rx_data) |=> (int_address == $past(addr_param[AW-1:0])));
assert_a37: assert property(@(posedge clock) $rose(reset) |=> (int_address == 0));
assert_a38: assert property(@(posedge clock) disable iff (reset) (bin_write_op && !addr_auto_inc) |=> $stable(int_address));
assert_a39: assert property(@(posedge clock) reset |-> (int_address == 0));
assert_a40: assert property(@(posedge clock) disable iff (reset) !(reset || ((main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) || ((main_sm == `MAIN_BIN_LEN) && new_rx_data)) |=> $stable(int_address));
assert_a41: assert property(@(posedge clock) ((main_sm == `MAIN_BIN_LEN) && new_rx_data) |=> (int_address == addr_param[AW-1:0]));
assert_a42: assert property(@(posedge clock) $fell(int_read || int_write) |-> !int_gnt);
assert_a43: assert property(@(posedge clock) $stable(int_req) |-> $stable(int_gnt));
assert_a44: assert property(@(posedge clock) $fell(int_req) |=> !int_gnt);
assert_a45: assert property(@(posedge clock) disable iff (reset) int_req |-> ##[1:2] int_gnt);
assert_a46: assert property(@(posedge clock) (int_gnt && (int_read || int_write)) |-> ##[1:2] int_gnt);
assert_a47: assert property(@(posedge clock) (int_gnt && int_write && $changed(int_wr_data)) |-> ##[1:2] $stable(int_gnt));
assert_a48: assert property(@(posedge clock) (int_wr_data == 0) && !int_req |-> !int_gnt);
assert_a49: assert property(@(posedge clock) disable iff (reset) int_req |-> ##[1:3] int_gnt);
assert_a50: assert property(@(posedge clock) int_req |-> int_gnt[*1:8]);
assert_a51: assert property(@(posedge clock) $changed(int_address) |-> !int_gnt);
assert_a52: assert property(@(posedge clock) int_gnt |-> (int_req && (int_read || int_write)));
assert_a53: assert property(@(posedge clock) !(reset && int_gnt));
assert_a54: assert property(@(posedge clock) $fell(reset) |=> !int_gnt);
assert_a55: assert property(@(posedge clock) reset |-> !int_gnt);
assert_a56: assert property(@(posedge clock) disable iff (reset) (int_req && !reset) |-> ##[1:4] int_gnt);
assert_a57: assert property(@(posedge clock) $fell(int_req) |-> ##[0:1] !int_gnt);
assert_a58: assert property(@(posedge clock) (int_gnt && $changed(int_address)) |=> int_gnt);
assert_a59: assert property(@(posedge clock) disable iff (reset) (int_req && !reset) |-> ##[1:3] int_gnt);
assert_a60: assert property(@(posedge clock) disable iff (!reset) !(reset && int_gnt));
assert_a61: assert property(@(posedge clock) int_gnt |-> (int_write || int_read));
assert_a62: assert property(@(posedge clock) disable iff (reset) $fell(int_req) |-> ##1 !int_gnt);
assert_a63: assert property(@(posedge clock) disable iff (reset) int_gnt |-> ##[0:7] !int_gnt);
assert_a64: assert property(@(posedge clock) disable iff (reset) ($rose(int_req) ##1 int_req[*4]) |-> (int_gnt [*1:5]));
assert_a65: assert property(@(posedge clock) disable iff (reset) (int_gnt && int_read) |-> ##[1:3] $stable(int_rd_data));
assert_a66: assert property(@(posedge clock) disable iff (reset) $fell(int_req) |-> ##[1:2] $fell(int_gnt));
assert_a67: assert property(@(posedge clock) $rose(reset) |-> ##1 !int_gnt);
assert_a68: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt) |-> int_gnt throughout int_read[->1]);
assert_a69: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt) |-> (int_rd_data >= 8'h00 && int_rd_data <= 8'hFF));
assert_a70: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt && (int_rd_data == 0)) |=> (int_rd_data != 0));
assert_a71: assert property(@(posedge clock) disable iff (reset) $fell(reset) |-> (int_rd_data == 0) until (int_read && int_gnt));
assert_a72: assert property(@(posedge clock) disable iff (reset) $fell(reset) |-> ##3 (int_rd_data >= 0 && int_rd_data <= 63));
assert_a73: assert property(@(posedge clock) disable iff (reset) !int_gnt |-> $stable(int_rd_data));
assert_a74: assert property(@(posedge clock) disable iff (reset) $changed(int_rd_data) |-> (int_read && int_gnt));
assert_a75: assert property(@(posedge clock) disable iff (reset) $fell(int_gnt) |-> $stable(int_rd_data)[*1]);
assert_a76: assert property(@(posedge clock) disable iff (reset) (int_gnt && $past(int_read) && int_read) |-> !$isunknown(int_rd_data));
assert_a77: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt) |-> $changed(int_rd_data));
assert_a78: assert property(@(posedge clock) disable iff (reset) $changed(int_rd_data) |-> $past(int_gnt));
assert_a79: assert property(@(posedge clock) disable iff (reset) int_read && int_gnt |=> $stable(int_rd_data)[*1]);
assert_a80: assert property(@(posedge clock) disable iff (reset) !int_read |-> $stable(int_rd_data));
assert_a81: assert property(@(posedge clock) disable iff (reset) int_read && !int_gnt |-> $stable(int_rd_data));
assert_a82: assert property(@(posedge clock) disable iff (reset) (!int_read || !int_gnt) && ($changed(ser_in) || $changed(ser_out)) |-> $stable(int_rd_data));
assert_a83: assert property(@(posedge clock) reset |-> (int_rd_data == 0));
assert_a84: assert property(@(posedge clock) disable iff (reset) $fell(int_read && int_gnt) |-> $stable(int_rd_data)[*1]);
assert_a85: assert property(@(posedge clock) disable iff (reset) ($rose(int_read) && int_gnt) |=> $stable(int_rd_data)[*1]);
assert_a86: assert property(@(posedge clock) reset |-> $stable(int_rd_data));
assert_a87: assert property(@(posedge clock) disable iff (reset) int_write |-> $stable(int_rd_data));
assert_a88: assert property(@(posedge clock) disable iff (reset) !int_gnt |-> int_rd_data === 8'bz);
assert_a89: assert property(@(posedge clock) disable iff (reset) !int_read && $changed(int_address) |-> $stable(int_rd_data));
assert_a90: assert property(@(posedge clock) disable iff (reset) $changed(int_rd_data) |-> $past(int_read && int_gnt));
assert_a91: assert property(@(posedge clock) $rose(!reset) |-> (int_rd_data == 0));
assert_a92: assert property(@(posedge clock) disable iff (reset) $fell(int_read) |-> $stable(int_rd_data)[*1]);
assert_a93: assert property(@(posedge clock) disable iff (reset) $fell(int_gnt) |-> $stable(int_rd_data)[*2]);
assert_a94: assert property(@(posedge clock) disable iff (reset) (!int_read || !int_gnt) && $changed(int_address) |-> $stable(int_rd_data));
assert_a95: assert property(@(posedge clock) disable iff (reset) $fell(int_req) && int_gnt |-> $stable(int_rd_data));
assert_a96: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt) |-> ##[1:2] $changed(int_rd_data));
assert_a97: assert property(@(posedge clock) disable iff (reset) !reset |-> (int_rd_data >= 0 && int_rd_data <= 255));
assert_a98: assert property(@(posedge clock) reset |-> ##1 (int_rd_data == 0));
assert_a99: assert property(@(posedge clock) (int_read && int_gnt) |-> ##[1:2] $changed(int_rd_data));
assert_a100: assert property(@(posedge clock) $changed(int_rd_data) |-> (int_read && int_gnt && !reset));
assert_a101: assert property(@(posedge clock) $rose(reset) |-> $stable(int_rd_data));
assert_a102: assert property(@(posedge clock) (!int_read && !int_write) |-> int_rd_data === 'z);
assert_a103: assert property(@(posedge clock) !(int_read && int_gnt) |-> int_rd_data === 'z);
assert_a104: assert property(@(posedge clock) int_rd_data !== 'z |-> (int_gnt && int_read));
assert_a105: assert property(@(posedge clock) (int_read && int_gnt) |=> (int_rd_data >= 0 && int_rd_data <= 255));
assert_a106: assert property(@(posedge clock) $changed(int_write) && !int_read |-> $stable(int_rd_data));
assert_a107: assert property(@(posedge clock) (int_rd_data >= 128 && int_rd_data <= 255) |=> (int_rd_data >= 64 && int_rd_data <= 255));
assert_a108: assert property(@(posedge clock) int_write |-> $stable(int_rd_data));
assert_a109: assert property(@(posedge clock) $fell(int_gnt) && int_read |=> $stable(int_rd_data));
assert_a110: assert property(@(posedge clock) (int_read && int_gnt) && $changed(ser_out) |-> $stable(int_rd_data));
assert_a111: assert property(@(posedge clock) $fell(int_read) |-> $past(int_rd_data) === int_rd_data);
assert_a112: assert property(@(posedge clock) int_read && $fell(int_req) && !int_gnt |-> $stable(int_rd_data));
assert_a113: assert property(@(posedge clock) ($rose(int_gnt) && int_read) |-> ##[1:3] (int_rd_data != 0));
assert_a114: assert property(@(posedge clock) $rose(!reset) |-> (int_rd_data === 8'b0));
assert_a115: assert property(@(posedge clock) int_read && !int_gnt |-> $stable(int_rd_data));
assert_a116: assert property(@(posedge clock) $changed(ser_out) |-> $stable(int_rd_data));
assert_a117: assert property(@(posedge clock) int_gnt && int_read |-> $stable(int_rd_data));
assert_a118: assert property(@(posedge clock) int_gnt && $changed(int_read) |-> $stable(int_rd_data));
assert_a119: assert property(@(posedge clock) (int_read && int_gnt && $fell(int_req)) |-> $changed(int_rd_data) [->1]);
assert_a120: assert property(@(posedge clock) (int_rd_data !== 'z) <-> (int_read && int_gnt));
assert_a121: assert property(@(posedge clock) (int_read && int_gnt) |-> $changed(int_rd_data) [->1]);
assert_a122: assert property(@(posedge clock) $changed(int_wr_data) && !int_write |-> $stable(int_rd_data));
assert_a123: assert property(@(posedge clock) (int_read && int_gnt) && $changed(int_address) |-> $stable(int_rd_data));
assert_a124: assert property(@(posedge clock) (int_read && int_gnt) && $changed(int_wr_data) |-> $stable(int_rd_data));
assert_a125: assert property(@(posedge clock) $changed(ser_in) && !(int_read && int_gnt) |-> $stable(int_rd_data));
assert_a126: assert property(@(posedge clock) disable iff (reset) $rose(int_write) && !int_read |-> $stable(int_rd_data));
assert_a127: assert property(@(posedge clock) disable iff (reset) (int_req && !int_gnt) |=> $stable(int_rd_data));
assert_a128: assert property(@(posedge clock) reset |-> !$isunknown(int_rd_data) && int_rd_data == 0);
assert_a129: assert property(@(posedge clock) disable iff (reset) $fell(int_gnt) |=> $stable(int_rd_data));
assert_a130: assert property(@(posedge clock) disable iff (reset) int_req && !int_gnt |-> $stable(int_rd_data));
assert_a131: assert property(@(posedge clock) disable iff (reset) $changed(int_req) && !int_gnt |-> $stable(int_rd_data));
assert_a132: assert property(@(posedge clock) disable iff (reset) $fell(int_gnt) && $past(int_read) |-> $stable(int_rd_data));
assert_a133: assert property(@(posedge clock) disable iff (reset) !int_gnt |-> !$isunknown(int_rd_data) && $stable(int_rd_data));
assert_a134: assert property(@(posedge clock) disable iff (reset) $changed(int_wr_data) && !int_read |-> $stable(int_rd_data));
assert_a135: assert property(@(posedge clock) disable iff (reset) !int_read && !int_gnt |-> $stable(int_rd_data));
assert_a136: assert property(@(posedge clock) disable iff (reset) $fell(int_read) && int_gnt |-> $stable(int_rd_data));
assert_a137: assert property(@(posedge clock) disable iff (reset) $changed(int_wr_data) && !int_write |-> $stable(int_rd_data));
assert_a138: assert property(@(posedge clock) disable iff (reset) !int_read && !int_gnt && $changed(ser_out) |-> $stable(int_rd_data));
assert_a139: assert property(@(posedge clock) disable iff (reset) $changed(ser_in) && !(int_read && int_gnt) |-> $stable(int_rd_data));
assert_a140: assert property(@(posedge clock) disable iff (reset) !$past(int_read) |-> int_rd_data == 0);
assert_a141: assert property(@(posedge clock) disable iff (reset) $fell(int_read) |=> $stable(int_rd_data));
assert_a142: assert property(@(posedge clock) disable iff (reset) int_read && int_gnt && $changed(ser_out) |-> $stable(int_rd_data));
assert_a143: assert property(@(posedge clock) disable iff (reset) (int_rd_data >= 0 && int_rd_data <= 127) |=> (int_rd_data >= 0 && int_rd_data <= 255));
assert_a144: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt) |-> int_rd_data == expected_data(int_address));
assert_a145: assert property(@(posedge clock) disable iff (reset) int_gnt && $fell(int_read) |-> $stable(int_rd_data));
assert_a146: assert property(@(posedge clock) disable iff (reset) $rose(int_read && int_gnt) |=> $changed(int_rd_data));
assert_a147: assert property(@(posedge clock) disable iff (reset) $fell(int_read) |-> ##[0:2] $stable(int_rd_data));
assert_a148: assert property(@(posedge clock) disable iff (reset) $changed(int_address) && !(int_read && int_gnt) |-> $stable(int_rd_data));
assert_a149: assert property(@(posedge clock) disable iff (reset) int_read && int_gnt |=> $stable(int_rd_data)[*1:$] until $fell(int_read));
assert_a150: assert property(@(posedge clock) $fell(reset) |-> ##2 (int_rd_data >= 0 && int_rd_data <= 255));
assert_a151: assert property(@(posedge clock) reset |=> int_rd_data == 0);
assert_a152: assert property(@(posedge clock) disable iff (reset) $changed(int_req) && !int_gnt |=> $stable(int_rd_data));
assert_a153: assert property(@(posedge clock) disable iff (reset) int_req && !int_gnt |-> !$isunknown(int_rd_data));
assert_a154: assert property(@(posedge clock) disable iff (reset) !int_gnt |-> !$isunknown(int_rd_data));
assert_a155: assert property(@(posedge clock) disable iff (reset) $rose(int_read && int_gnt) |-> ##[1:2] $changed(int_rd_data));
assert_a156: assert property(@(posedge clock) reset |-> int_rd_data == 0);
assert_a157: assert property(@(posedge clock) (int_read && !int_req) |=> !int_read);
assert_a158: assert property(@(posedge clock) int_read |=> !int_read);
assert_a159: assert property(@(posedge clock) (int_read && int_req && int_gnt) |=> !int_read);
assert_a160: assert property(@(posedge clock) int_read |=> $past(int_rd_data,1) == $past(int_rd_data,2));
assert_a161: assert property(@(posedge clock) int_read |-> !$isunknown(int_address));
assert_a162: assert property(@(posedge clock) !int_req |-> !int_read);
assert_a163: assert property(@(posedge clock) int_read |-> $past(int_address,1) == int_address);
assert_a164: assert property(@(posedge clock) int_read |=> $stable(int_rd_data));
assert_a165: assert property(@(posedge clock) $stable(int_gnt) && int_gnt |-> !int_read);
assert_a166: assert property(@(posedge clock) (int_read && int_req && int_gnt) |=> !int_read);
assert_a167: assert property(@(posedge clock) (int_read && int_req && int_gnt) |=> !int_read throughout !(int_req && int_gnt)[->1]);
assert_a168: assert property(@(posedge clock) reset |-> !int_read);
assert_a169: assert property(@(posedge clock) !(int_read && int_write));
assert_a170: assert property(@(posedge clock) int_read |-> $stable(int_address));
assert_a171: assert property(@(posedge clock) (int_read && $stable(int_address)) |=> !(int_read && $stable(int_address)));
assert_a172: assert property(@(posedge clock) int_read |-> (int_req && int_gnt));
assert_a173: assert property(@(posedge clock) $rose(int_read) |-> $stable(int_address)[*1]);
assert_a174: assert property(@(posedge clock) $rose(int_read) |-> (int_req throughout ( ##[0:$] $fell(int_req) )));
assert_a175: assert property(@(posedge clock) $stable(int_gnt) && int_gnt |-> !int_read);
assert_a176: assert property(@(posedge clock) $rose(int_read) |-> $past(int_req));
assert_a177: assert property(@(posedge clock) $rose(int_read) |-> (int_req && int_gnt));
assert_a178: assert property(@(posedge clock) !(int_read && int_write));
assert_a179: assert property(@(posedge clock) reset |-> !int_read);
assert_a180: assert property(@(posedge clock) int_read |-> int_gnt);
assert_a181: assert property(@(posedge clock) int_read |-> (int_req && int_gnt));
assert_a182: assert property(@(posedge clock) disable iff (reset) ($rose(int_req) && !int_gnt [*5]) |-> ##1 !int_req);
assert_a183: assert property(@(posedge clock) disable iff (reset) (int_req && (int_write || int_read)) |-> !int_gnt until !(int_write || int_read));
assert_a184: assert property(@(posedge clock) (int_req && (int_read || int_write)) |-> int_gnt);
assert_a185: assert property(@(posedge clock) $rose(int_req) |-> ##1 int_req);
assert_a186: assert property(@(posedge clock) int_req |-> !int_gnt);
assert_a187: assert property(@(posedge clock) disable iff (reset) ($fell(int_gnt)) |-> ##[0:2] !int_req);
assert_a188: assert property(@(posedge clock) disable iff (reset) (int_req && !int_gnt) |-> ##1 !int_req);
assert_a189: assert property(@(posedge clock) disable iff (reset) (int_req && int_gnt) |-> (int_rd_data == int_address || int_wr_data == int_address));
assert_a190: assert property(@(posedge clock) !(int_req && int_write));
assert_a191: assert property(@(posedge clock) int_req |-> (int_read || int_write));
assert_a192: assert property(@(posedge clock) disable iff (reset) int_rd_data |-> !int_req);
assert_a193: assert property(@(posedge clock) disable iff (reset) (int_rd_data || int_wr_data) |-> !int_req);
assert_a194: assert property(@(posedge clock) $rose(reset) |-> !int_req);
assert_a195: assert property(@(posedge clock) disable iff (reset) int_req |-> (int_address != 0));
assert_a196: assert property(@(posedge clock) $rose(!reset) |=> !int_req[*2]);
assert_a197: assert property(@(posedge clock) disable iff (reset) int_req |-> ##[1:3] int_gnt);
assert_a198: assert property(@(posedge clock) disable iff (reset) ((int_rd_data && !int_read) || (int_wr_data && !int_write)) |-> !int_req);
assert_a199: assert property(@(posedge clock) reset |-> !int_req);
// assert_a200: assert property(@(posedge clock) disable iff (reset) $rose(int_req) |-> ($stable(int_address) throughout (int_req until int_gnt)));
assert_a201: assert property(@(posedge clock) $fell(reset) |-> ##2 !int_req);
assert_a202: assert property(@(posedge clock) disable iff (reset) $fell(int_req) |-> ##1 !int_gnt);
assert_a203: assert property(@(posedge clock) disable iff (reset) (int_req && ser_in) |-> ##[1:2] int_gnt);
assert_a204: assert property(@(posedge clock) $rose(reset) |-> ##1 !int_req);
assert_a205: assert property(@(posedge clock) disable iff (reset) (int_req && int_read) |-> ##[1:3] int_gnt);
assert_a206: assert property(@(posedge clock) disable iff (reset) int_req |=> (int_req throughout int_gnt[->1]) or reset);
assert_a207: assert property(@(posedge clock) disable iff (reset) (int_req && !int_gnt) |-> $stable(int_wr_data) throughout (int_req[*1:$] ##0 int_gnt));
assert_a208: assert property(@(posedge clock) disable iff (reset) !write_req && !reset |=> $stable(int_wr_data));
assert_a209: assert property(@(posedge clock) disable iff (reset) $changed(int_wr_data) |=> ##1 $stable(int_wr_data) or reset);
assert_a210: assert property(@(posedge clock) disable iff (reset) (write_op || bin_write_op) && !new_rx_data |=> $stable(int_wr_data));
assert_a211: assert property(@(posedge clock) disable iff (reset) (write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) |=> (int_wr_data == $past(data_param)));
assert_a212: assert property(@(posedge clock) disable iff (reset) write_op && !data_in_hex_range && !bin_write_op |=> (int_wr_data == $past(data_param)));
assert_a213: assert property(@(posedge clock) reset |-> (int_wr_data == 0) [*1:$] until !reset);
assert_a214: assert property(@(posedge clock) disable iff (reset) (bin_write_op && (main_sm == `MAIN_BIN_DATA) && new_rx_data) |=> (int_wr_data == $past(rx_data)));
assert_a215: assert property(@(posedge clock) disable iff (reset) $changed(int_wr_data) |-> ##[1:$] $stable(int_wr_data)[*1]);
assert_a216: assert property(@(posedge clock) disable iff (reset) new_rx_data && !(main_sm == `MAIN_ADDR || main_sm == `MAIN_BIN_DATA) |=> $stable(int_wr_data));
assert_a217: assert property(@(posedge clock) disable iff (reset) (write_op || bin_write_op) |=> $changed(int_wr_data));
assert_a218: assert property(@(posedge clock) disable iff (reset) write_op && !new_rx_data |=> $stable(int_wr_data));
assert_a219: assert property(@(posedge clock) disable iff (reset) !(write_op || bin_write_op) && (main_sm == `MAIN_ADDR || main_sm == `MAIN_BIN_DATA) |=> $stable(int_wr_data));
assert_a220: assert property(@(posedge clock) disable iff (reset) ($rose(write_op)) ##1 (write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) |=> (int_wr_data == $past(data_param)));
assert_a221: assert property(@(posedge clock) reset |=> (int_wr_data == 0) and (!reset throughout (write_op || bin_write_op)[->1]) |=> $stable(int_wr_data));
assert_a222: assert property(@(posedge clock) disable iff (reset) !reset && !(write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) && !(bin_write_op && (main_sm == `MAIN_BIN_DATA) && new_rx_data) |=> ($stable(int_wr_data)));
assert_a223: assert property(@(posedge clock) disable iff (reset) ($changed(int_wr_data)) |=> ($stable(int_wr_data)[*1] or (write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) or (bin_write_op && (main_sm == `MAIN_BIN_DATA) && new_rx_data)));
assert_a224: assert property(@(posedge clock) disable iff (reset) (write_op && (main_sm != `MAIN_ADDR)) |=> ($stable(int_wr_data)));
assert_a225: assert property(@(posedge clock) disable iff (reset) ($fell(write_req)) |-> ##[1:2] ($stable(int_wr_data)));
assert_a226: assert property(@(posedge clock) disable iff (reset) ($changed(write_op) || $changed(bin_write_op)) |-> $stable(int_wr_data));
assert_a227: assert property(@(posedge clock) disable iff (reset) $rose(write_op || bin_write_op) |-> !$isunknown(int_wr_data));
assert_a228: assert property(@(posedge clock) reset |-> (int_wr_data == 0));
assert_a229: assert property(@(posedge clock) $changed(int_wr_data) |-> $past(write_op || bin_write_op));
assert_a230: assert property(@(posedge clock) disable iff (reset) $changed(int_wr_data) |-> ($past(new_rx_data) && ($past(write_op) || $past(bin_write_op))));
assert_a231: assert property(@(posedge clock) $rose(!reset) |=> (int_wr_data == 0) until $rose(write_op));
assert_a232: assert property(@(posedge clock) disable iff (reset) $changed(int_wr_data) |-> ($past(write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) || $past(bin_write_op && (main_sm == `MAIN_BIN_DATA) && new_rx_data)));
assert_a233: assert property(@(posedge clock) (write_op && bin_write_op) |-> if (main_sm == `MAIN_ADDR) (int_wr_data == data_param) else if (main_sm == `MAIN_BIN_DATA) (int_wr_data == rx_data));
assert_a234: assert property(@(posedge clock) disable iff (reset) !(write_op || bin_write_op) |=> $stable(int_wr_data));
assert_a235: assert property(@(posedge clock) (write_op && (main_sm == `MAIN_ADDR) && new_rx_data && !data_in_hex_range) |=> (int_wr_data == $past(data_param)));
assert_a236: assert property(@(posedge clock) reset |=> (int_wr_data == 0));
assert_a237: assert property(@(posedge clock) disable iff (reset) (bin_write_op && (main_sm != `MAIN_BIN_DATA)) |=> $stable(int_wr_data));
assert_a238: assert property(@(posedge clock) $fell(reset) |=> (int_wr_data == 0) until (write_op || bin_write_op));
assert_a239: assert property(@(posedge clock) (int_gnt && write_req) |=> int_write);
assert_a240: assert property(@(posedge clock) (int_gnt && write_req) |-> (int_write && !write_req));
assert_a241: assert property(@(posedge clock) (int_gnt && write_req) |=> int_write ##1 !int_write);
assert_a242: assert property(@(posedge clock) (!write_req && int_gnt) |=> !int_write);
assert_a243: assert property(@(posedge clock) (int_write && !write_req) |=> !int_write);
assert_a244: assert property(@(posedge clock) $stable(int_gnt) && $stable(write_req) |-> $stable(int_write));
assert_a245: assert property(@(posedge clock) (!int_gnt && !write_req) |=> !int_write);
assert_a246: assert property(@(posedge clock) reset |=> !int_write);
assert_a247: assert property(@(posedge clock) (int_gnt && write_req) |=> (int_write && !write_req));
assert_a248: assert property(@(posedge clock) (int_write && !(int_gnt && write_req)) |=> !int_write);
assert_a249: assert property(@(posedge clock) !write_req |-> !int_write);
assert_a250: assert property(@(posedge clock) $rose(int_gnt) && !write_req |-> !int_write);
assert_a251: assert property(@(posedge clock) $fell(int_gnt) && write_req |=> !int_write);
assert_a252: assert property(@(posedge clock) int_write |-> int_gnt && write_req);
assert_a253: assert property(@(posedge clock) int_write |=> (int_gnt && write_req) || !int_write);
assert_a254: assert property(@(posedge clock) int_gnt && !write_req |=> !int_write);
assert_a255: assert property(@(posedge clock) reset |-> !int_write);
assert_a256: assert property(@(posedge clock) write_req && !int_gnt |=> !int_write);
assert_a257: assert property(@(posedge clock) disable iff (reset) int_write == (int_gnt && write_req));
assert_a258: assert property(@(posedge clock) disable iff (reset) (!int_gnt || !write_req) |=> !int_write);
assert_a259: assert property(@(posedge clock) $rose(!reset) |=> (int_write == (int_gnt && write_req)));
assert_a260: assert property(@(posedge clock) disable iff (reset) (int_gnt && write_req) |=> (int_write && !write_req));
assert_a261: assert property(@(posedge clock) disable iff (reset) (!int_gnt && write_req) |=> !int_write);
assert_a262: assert property(@(posedge clock) disable iff (reset) (bin_write_op && (main_sm == MAIN_BIN_DATA) && new_rx_data) |=> write_req);
assert_a263: assert property(@(posedge clock) (reset && int_gnt && write_req) |=> !int_write);
assert_a264: assert property(@(posedge clock) $rose(reset) |=> (rx_data == 8'h0));
assert_a265: assert property(@(posedge clock) $fell(reset) |=> $stable(ser_out)[*2]);
assert_a266: assert property(@(posedge clock) $fell(reset) ##1 (rx_busy && ce_1_mid) |=> (data_buf != $past(data_buf)));
assert_a267: assert property(@(posedge clock) reset |-> !int_gnt);
assert_a268: assert property(@(posedge clock) reset throughout (##[1:$] !reset) |-> $stable(rx_data));
assert_a269: assert property(@(posedge clock) $rose(reset) |=> (!int_write && !int_read));
assert_a270: assert property(@(posedge clock) $rose(reset) |=> !tx_busy);
assert_a271: assert property(@(posedge clock) $rose(reset) |=> (new_rx_data == 1'b0));
assert_a272: assert property(@(posedge clock) reset |-> !(rx_busy && ce_1_mid && !reset));
assert_a273: assert property(@(posedge clock) $rose(reset) |=> (int_rd_data == '0));
assert_a274: assert property(@(posedge clock) $rose(reset) |=> (int_address == '0));
assert_a275: assert property(@(posedge clock) disable iff (reset) !new_rx_data throughout (1'b1)[*0:$] until (valid_reception_condition));
// assert_a276: assert property(@(posedge clock) $rose(reset) |-> (rx_data == 8'h0 && new_rx_data == 1'b0 && data_buf == 8'h0) regardless_of (ser_in));
assert_a277: assert property(@(posedge clock) $fell(reset) |=> $stable(rx_data) until (rx_data_change_condition));
assert_a278: assert property(@(posedge clock) $rose(reset) |=> (rx_data == 8'h0 && new_rx_data == 1'b0 && data_buf == 8'h0));
assert_a279: assert property(@(posedge clock) $rose(reset) |=> !int_req);
assert_a280: assert property(@(posedge clock) $fell(reset) |-> ##[1:3] $changed(ser_in));
assert_a281: assert property(@(posedge clock) reset |-> (!int_write && !int_read));
assert_a282: assert property(@(posedge clock) $rose(reset) |=> (data_buf == 8'h0));
assert_a283: assert property(@(posedge clock) $rose(reset) |-> reset[*2]);
assert_a284: assert property(@(posedge clock) $fell(reset) |=> $stable(rx_data) && $stable(data_buf));
assert_a285: assert property(@(posedge clock) $rose(reset) |=> !new_rx_data);
assert_a286: assert property(@(posedge clock) $rose(reset) |=> (int_rd_data == 8'h0));
assert_a287: assert property(@(posedge clock) $rose(reset) |=> $stable(ser_out) throughout (reset[*1:$]));
// assert_a288: assert property(@(posedge clock) disable iff (reset) $rose(ser_in) && $fell(ser_in) within [0:$] |-> $stable(ser_out));
assert_a289: assert property(@(posedge clock) disable iff (reset) (!tx_busy) |-> ##4 (ser_out == $past(ser_in,4)));
assert_a290: assert property(@(posedge clock) disable iff (reset || !ce_16) ($fell(ser_in) ##1 !$rose(ser_in)[*10]) |-> !new_rx_data);
assert_a291: assert property(@(posedge clock) disable iff (reset) $fell(ser_in) |-> ##[1:16] int_req);
// assert_a292: assert property(@(posedge clock) disable iff (reset) ($rose(ser_in) && $fell(ser_in) within [0:$]) |-> $stable(int_wr_data));
assert_a293: assert property(@(posedge clock) disable iff (reset) (ser_in == 0)[*16] |-> $stable(int_address));
// assert_a294: assert property(@(posedge clock) disable iff (reset) ($stable(ser_in)[*8] && int_req) |-> ##1 int_gnt);
assert_a295: assert property(@(posedge clock) (reset) |-> $stable(ser_in));
assert_a296: assert property(@(posedge clock) disable iff (reset) ($fell(ser_in) ##1 $changed(ser_in)[*8]) |-> ##[1:16] int_write);
// assert_a297: assert property(@(posedge ce_16) $rose(ser_in) && $fell(ser_in) within [0:$] |-> $stable(ser_in));
// assert_a298: assert property(@(posedge clock) $rose(!reset) |-> $stable(ser_in, 2));
assert_a299: assert property(@(posedge clock) reset |-> (ser_out == $past(ser_out,1)) and (!$changed(int_write)) and (!$changed(int_read)));
assert_a300: assert property(@(posedge clock) disable iff (reset) (int_read && $fell(ser_in)) |=> (int_read throughout !$fell(ser_in))[*1:$] ##1 $fell(ser_in));
assert_a301: assert property(@(posedge clock) disable iff (reset) ser_in[*10] |-> !int_read);
assert_a302: assert property(@(posedge clock) disable iff (reset) $fell(ser_in) |-> ##[1:3] int_req);
assert_a303: assert property(@(posedge clock) disable iff (reset) (ser_in == 0) throughout (ce_16[->24]) |-> framing_error);
// assert_a304: assert property(@(posedge clock) disable iff (reset) $rose(!reset) ##4 (!reset throughout (($stable(ser_in, 2)) or ($fell(ser_in) ##2 $stable(ser_in)))));
assert_a305: assert property(@(posedge clock) disable iff (reset) $fell(ser_in) ##[1:$] $rose(ser_in) |-> ##[0:16] int_write [*1] ##1 !int_write);
assert_a306: assert property(@(posedge clock) ($fell(reset) && (ser_in == 0)) ##1 (ser_in == 1)[*4] |-> !framing_error);
assert_a307: assert property(@(posedge clock) disable iff (reset) (frame_end && ce_16) |-> ##[1:2] new_rx_data);
assert_a308: assert property(@(posedge clock) $rose(!reset) |-> strong(##[0:16] $stable(ser_in)));
assert_a309: assert property(@(posedge clock) disable iff (reset) ($fell(ser_in) ##1 ser_in[*8]) |-> ##[1:24] (int_wr_data == $past(ser_in, 8)));
assert_a310: assert property(@(posedge clock) disable iff (reset) $fell(ser_in) && ce_16 |-> ##[1:16] $rose(ser_in));
assert_a311: assert property(@(posedge clock) disable iff (reset) $fell(ser_in) |-> ##[1:16] (new_rx_data && $stable(ser_out)));
assert_a312: assert property(@(posedge clock) disable iff (reset) ($countones(ser_in) >= 10) |-> $stable(ser_in) until $fell(ser_in));
assert_a313: assert property(@(posedge clock) disable iff (reset) ($countones(ser_in) >= 16) |-> ##[1:16] !int_read);
// assert_a314: assert property(@(posedge clock) disable iff (reset) (ser_in == 1'b0 ##1 ser_in == 1'b1 ##1 ser_in == 1'b0 ##1 ser_in == 1'b1 ##1 ser_in == 1'b0 ##1 ser_in == 1'b1 ##1 ser_in == 1'b0 ##1 ser_in == 1'b1) && ce_16 |-> (int_address == 8'h55));
assert_a315: assert property(@(posedge clock) reset |-> $stable(int_rd_data));
assert_a316: assert property(@(posedge clock) disable iff (reset) ($fell(ser_in) && ce_16) |-> ##[1:$] (new_rx_data && $stable(ce_16)[*1:$]));
assert_a317: assert property(@(posedge clock) disable iff (reset) ($rose(ser_in) && int_req) |-> ##[1:2] !int_gnt);
assert_a318: assert property(@(posedge clock) $rose(int_gnt) |-> ##[1:2] $stable(ser_out));
assert_a319: assert property(@(posedge clock) int_write |-> ##[1:2] (ser_out == 0 || ser_out == 1));
assert_a320: assert property(@(posedge clock) int_gnt && !int_req |-> $stable(ser_out));
assert_a321: assert property(@(posedge clock) (int_req && !int_gnt) |-> ##5 ($stable(ser_out)[*5]));
assert_a322: assert property(@(posedge clock) (int_req && !int_gnt) |-> ##[1:10] $changed(ser_out));
assert_a323: assert property(@(posedge clock) reset |-> $stable(ser_out));
assert_a324: assert property(@(posedge clock) (int_read && int_write) |-> $stable(ser_out));
assert_a325: assert property(@(posedge clock) $fell(reset) |-> (ser_out == 0)[*3]);
assert_a326: assert property(@(posedge clock) (!int_read && !int_write) |-> ##4 ($fell(ser_out) || $rose(ser_out))[*4]);
assert_a327: assert property(@(posedge clock) $changed(int_address) && !int_write |-> $stable(ser_out));
assert_a328: assert property(@(posedge clock) $changed(int_read) || $changed(int_write) |-> ##1 !$isunknown(ser_out) throughout ##[0:1] $stable(ser_out));
assert_a329: assert property(@(posedge clock) disable iff (reset) $changed(ser_out) |-> $rose(clock));
assert_a330: assert property(@(posedge clock) (int_req && !int_gnt) |-> $stable(ser_out));
assert_a331: assert property(@(posedge clock) int_write |-> ser_out == int_wr_data[0]);
assert_a332: assert property(@(posedge clock) reset |=> $stable(ser_out));
assert_a333: assert property(@(posedge clock) $fell(reset) |-> (ser_out == 1'b0));
assert_a334: assert property(@(posedge clock) $fell(int_write) |=> (ser_out == 1'b1));
assert_a335: assert property(@(posedge clock) ($changed(int_address) && int_write) |-> (ser_out == 1'b1)[->1] ##1 ser_out != 1'b1);
assert_a336: assert property(@(posedge clock) disable iff (int_write) (ser_in |-> ##1 ser_out == $past(ser_in)));
assert_a337: assert property(@(posedge clock) (int_req && int_gnt) |-> ##[1:4] !$stable(ser_out));
assert_a338: assert property(@(posedge clock) $rose(int_read) |-> ##[1:10] $changed(ser_out));
assert_a339: assert property(@(posedge clock) disable iff (reset) $changed(int_rd_data) |-> ##[1:2] $stable(ser_out));
assert_a340: assert property(@(posedge clock) disable iff (reset) int_write |-> (ser_out == int_wr_data[0]));
assert_a341: assert property(@(posedge clock) $fell(reset) |-> ##[1:2] (ser_out == 1'b1));
assert_a342: assert property(@(posedge clock) $rose(reset) |-> ##[0:2] ($stable(ser_out)) and $fell(reset) |-> ##[0:2] ($stable(ser_out)));
// assert_a343: assert property(@(posedge clock) disable iff (reset) (int_read && $changed(int_rd_data)) |-> ##[1:4] (ser_out == $past(int_rd_data, 4)[7:0]));
assert_a344: assert property(@(posedge clock) disable iff (reset) (int_write && int_gnt)[*3] |-> (ser_out == int_wr_data[7:0]));
assert_a345: assert property(@(posedge clock) disable iff (reset) $fell(int_read) |-> (ser_out == 1'b1)[*3]);
assert_a346: assert property(@(posedge clock) disable iff (reset) (int_read && int_gnt) |-> ##[1:3] (ser_out == $past(ser_in, 3)));
assert_a347: assert property(@(posedge clock) disable iff (reset) ($past(int_address) == 8'h00 && int_address != 8'h00) |-> ##[1:5] (ser_out == 1'b1));
assert_a348: assert property(@(posedge clock) disable iff (reset) int_read |-> (ser_out == ^int_rd_data));


endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------

// File: baud_gen.sv
//---------------------------------------------------------------------------------------
// baud rate generator for uart 
//
// this module has been changed to receive the baud rate dividing counter from registers.
// the two registers should be calculated as follows:
// first register:
// 		baud_freq = 16*baud_rate / gcd(global_clock_freq, 16*baud_rate)
// second register:
// 		baud_limit = (global_clock_freq / gcd(global_clock_freq, 16*baud_rate)) - baud_freq 
//
//---------------------------------------------------------------------------------------

module baud_gen 
(
	clock, reset, 
	ce_16, baud_freq, baud_limit 
);
//---------------------------------------------------------------------------------------
// modules inputs and outputs 
input 			clock;		// global clock input 
input 			reset;		// global reset input 
output			ce_16;		// baud rate multiplyed by 16 
input	[11:0]	baud_freq;	// baud rate setting registers - see header description 
input	[15:0]	baud_limit;

// internal registers 
reg ce_16;
reg [15:0]	counter;
//---------------------------------------------------------------------------------------
// module implementation 
// baud divider counter  
always @ (posedge clock or posedge reset)
begin
	if (reset) 
		counter <= 16'b0;
	else if (counter >= baud_limit) 
		counter <= counter - baud_limit;
	else 
		counter <= counter + baud_freq;
end

// clock divider output 
always @ (posedge clock or posedge reset)
begin
	if (reset)
		ce_16 <= 1'b0;
	else if (counter >= baud_limit) 
		ce_16 <= 1'b1;
	else 
		ce_16 <= 1'b0;
end 

endmodule
//---------------------------------------------------------------------------------------
//						Th.. Th.. Th.. Thats all folks !!!
//---------------------------------------------------------------------------------------
